--------------------------------------------------------------------------------
-- HEIG-VD, Haute Ecole d'Ingenierie et de Gestion du canton de Vaud
-- Institut REDS, Reconfigurable & Embedded Digital Systems
--
-- File         : cpt_pos.vhd
--
-- Description  : 
--
-- Author       : L. Fournier
-- Date         : 28.01.2023
-- Version      : 1.0
--
-- Use          : SysLog2 labo : Acqu pos
--
--| Modifications |-------------------------------------------------------------
-- Version   Auteur      Date               Description
-- 1.0       LFR         21.04.2023         Empty version.
--------------------------------------------------------------------------------

--| Library |-------------------------------------------------------------------
library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;
--------------------------------------------------------------------------------

--| Entity |--------------------------------------------------------------------
entity cpt_pos is
    port(
        clock_i    : in  std_logic; -- system clock
        reset_i    : in  std_logic; -- asynchronous reset
        -- A completer
    );
end cpt_pos;
--------------------------------------------------------------------------------

--| Architecture |--------------------------------------------------------------
architecture rtl of cpt_pos is

    --| Signals |---------------------------------------------------------------
   
    ----------------------------------------------------------------------------

begin

    --| Outputs affectation |---------------------------------------------------

    ----------------------------------------------------------------------------

end rtl;
--------------------------------------------------------------------------------