--------------------------------------------------------------------------------
-- HEIG-VD, Haute Ecole d'Ingenierie et de Gestion du canton de Vaud
-- Institut REDS, Reconfigurable & Embedded Digital Systems
--
-- File         : mss_det_rot.vhd
--
-- Description  : 
--
-- Author       : L. Fournier
-- Date         : 28.01.2023
-- Version      : 1.0
--
-- Use          : SysLog2 labo : Acqu pos
--
--| Modifications |-------------------------------------------------------------
-- Version   Auteur      Date               Description
-- 1.0       LFR         21.04.2023         Empty version.
--------------------------------------------------------------------------------

--| Library |-------------------------------------------------------------------
library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;
--------------------------------------------------------------------------------

--| Entity |--------------------------------------------------------------------
entity mss_det_rot is
    port(
        clock_i   : in  std_logic;
        reset_i   : in  std_logic;
        -- A completer
    );
end mss_det_rot;
--------------------------------------------------------------------------------

--| Architecture |--------------------------------------------------------------
architecture fsm of mss_det_rot is

    --| Types |-----------------------------------------------------------------

    ----------------------------------------------------------------------------

    --| Signals |---------------------------------------------------------------

    ----------------------------------------------------------------------------

begin

    --| Outputs affectation |---------------------------------------------------

    ----------------------------------------------------------------------------

end fsm;
--------------------------------------------------------------------------------